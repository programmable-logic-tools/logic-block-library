/**
 * This module calculates the tick numbers for turning the
 * highside and lowside switches of a half-bridge on and off
 * from the turn-on and -off durations and the deadtimes.
 */
